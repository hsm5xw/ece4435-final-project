CONFIGURATION memory_stage_struct_config OF memory_stage IS
   FOR struct
   END FOR;
END memory_stage_struct_config;