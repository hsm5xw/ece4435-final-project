CONFIGURATION SimpleMux3_Behavior_config OF SimpleMux3 IS
   FOR Behavior
   END FOR;
END SimpleMux3_Behavior_config;