CONFIGURATION lab10_WriteBack_Stage_struct_config OF lab10_WriteBack_Stage IS
   FOR struct
   END FOR;
END lab10_WriteBack_Stage_struct_config;