CONFIGURATION SRAM_behavior_config OF SRAM IS
   FOR behavior
   END FOR;
END SRAM_behavior_config;