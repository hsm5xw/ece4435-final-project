CONFIGURATION SimpleMux4_Behavior_config OF SimpleMux4 IS
   FOR Behavior
   END FOR;
END SimpleMux4_Behavior_config;