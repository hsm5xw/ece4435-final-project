CONFIGURATION mini_ALU_struct_config OF mini_ALU IS
   FOR struct
   END FOR;
END mini_ALU_struct_config;