CONFIGURATION mini_Shifter_Behavior_config OF mini_Shifter IS
   FOR Behavior
   END FOR;
END mini_Shifter_Behavior_config;