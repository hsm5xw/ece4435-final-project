CONFIGURATION Decoder_Behavior_config OF Decoder IS
   FOR Behavior
   END FOR;
END Decoder_Behavior_config;