CONFIGURATION ALU_ROM_Behavior_config OF ALU_ROM IS
   FOR Behavior
   END FOR;
END ALU_ROM_Behavior_config;