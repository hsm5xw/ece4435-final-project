CONFIGURATION Reg_Behavior_config OF Reg IS
   FOR Behavior
   END FOR;
END Reg_Behavior_config;