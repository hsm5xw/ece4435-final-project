CONFIGURATION Processor_Behavior_config OF Processor IS
   FOR Behavior
   END FOR;
END Processor_Behavior_config;