CONFIGURATION MemoryArbiter_struct_config OF MemoryArbiter IS
   FOR struct
   END FOR;
END MemoryArbiter_struct_config;