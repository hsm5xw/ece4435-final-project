CONFIGURATION Decode_ROM_Behavior_config OF Decode_ROM IS
   FOR Behavior
   END FOR;
END Decode_ROM_Behavior_config;