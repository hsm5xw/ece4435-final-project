CONFIGURATION SimpleMux2_Behavior_config OF SimpleMux2 IS
   FOR Behavior
   END FOR;
END SimpleMux2_Behavior_config;